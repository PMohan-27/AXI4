module axi4_lite_slave #(parameter DATA_WIDTH = 32, ADDRESS_WIDTH = 32)(
    // Global
    input ACLK,
    input ARESETn,
    
);


endmodule
