module axi4_lite(

);


endmodule